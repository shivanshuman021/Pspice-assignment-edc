*************Example4***************
Vin 1 0 DC 10V;
Is 4 3 DC 2A;
R1 1 2 5;
R2 2 3 10;
R3 2 0 20;
R4 3 4 40;
R5 5 0 10;
Vx 4 5 DC 0V;
.TF V(2,4) Vin;
.END;