* C:\Users\boruto_uz\Desktop\edc\q1\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Fri Feb 19 17:54:26 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
