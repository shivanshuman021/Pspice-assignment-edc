**************QUES9**********************
VGS 1 0 DC 5V;
VDS 2 0 DC 5V;
M1 2 1 0 0 MOS1 W=5u L=1u;
.MODEL MOS1 NMOS VTO=0.7 KP=110V LAMBDA=0.4 PHI=0.7 GAMMA=0;
.DC VDS 0 5 0.2 VGS 1 5 1;
.PROBE;
.END;
