************Example3.CIR*************
Vs 1 0 DC 20V;
Is 0 4 DC 50mA;
R1 1 2 500;
R2 2 5 800;
R3 2 4 1KOHM;
R4 4 0 200;
Vx 3 0 DC 0V;
Vy 5 4 DC 0V;
.DC Vs LIST 5V 20V 30V Is 50ma 150mA 50mA;
.PRINT DC V(4) I(Vx) I(Vy);
.PLOT DC I(Vy);
.PROBE;
.END