* C:\Users\boruto_uz\Desktop\edc\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Wed Feb 17 08:51:33 2021



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
