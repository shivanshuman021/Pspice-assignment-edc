******************QUE8***********************
IB 0 1 DC 1mA;
VCE 2 0 DC 12V;
Q1 2 1 0 Q2N2222A;
.MODEL Q2N2222A NPN (IS=2.105E-16 BF=173 VA=83.3V CJE=29.6PF CJC=19.4PF TF 489.88PS TR=4.9NS);
.DC VCE 0 10V 0.02V IB 0 1mA 200uA;
.PROBE;
.END;
